wire dec_xcr2gpr     = (encoded & 32'hfff8707f) == 32'h1000002b;
wire dec_gpr2xcr     = (encoded & 32'hfff0787f) == 32'h1100002b;
wire dec_init        = (encoded & 32'hffffffff) == 32'h1110082b;
wire dec_rngseed     = (encoded & 32'hfff87fff) == 32'h800002b;
wire dec_rngsamp     = (encoded & 32'hfffff87f) == 32'h810082b;
wire dec_rngtest     = (encoded & 32'hfffff07f) == 32'h820002b;
wire dec_cmov_t      = (encoded & 32'hff08787f) == 32'h1800082b;
wire dec_cmov_f      = (encoded & 32'hff08787f) == 32'h1800002b;
wire dec_padd        = (encoded & 32'h1f08787f) == 32'h600002b;
wire dec_psub        = (encoded & 32'h1f08787f) == 32'h600082b;
wire dec_pmul_l      = (encoded & 32'h1f08787f) == 32'he00002b;
wire dec_pmul_h      = (encoded & 32'h1f08787f) == 32'he00082b;
wire dec_pclmul_l    = (encoded & 32'h1f08787f) == 32'he08002b;
wire dec_pclmul_h    = (encoded & 32'h1f08787f) == 32'he08082b;
wire dec_psll        = (encoded & 32'h1f08787f) == 32'h1600002b;
wire dec_psrl        = (encoded & 32'h1f08787f) == 32'h1600082b;
wire dec_prot        = (encoded & 32'h1f08787f) == 32'h1608082b;
wire dec_psll_i      = (encoded & 32'h1e08787f) == 32'h1e00002b;
wire dec_psrl_i      = (encoded & 32'h1e08787f) == 32'h1e00082b;
wire dec_prot_i      = (encoded & 32'h1e08787f) == 32'h1e08082b;
wire dec_sha3_xy     = (encoded & 32'h3e00707f) == 32'hc00002b;
wire dec_sha3_x1     = (encoded & 32'h3e00707f) == 32'h1400002b;
wire dec_sha3_x2     = (encoded & 32'h3e00707f) == 32'h2400002b;
wire dec_sha3_x4     = (encoded & 32'h3e00707f) == 32'h1c00002b;
wire dec_sha3_yx     = (encoded & 32'h3e00707f) == 32'h3400002b;
wire dec_aessub_enc  = (encoded & 32'hff08787f) == 32'h400002b;
wire dec_aessub_encrot = (encoded & 32'hff08787f) == 32'h400082b;
wire dec_aessub_dec  = (encoded & 32'hff08787f) == 32'h408002b;
wire dec_aessub_decrot = (encoded & 32'hff08787f) == 32'h408082b;
wire dec_aesmix_enc  = (encoded & 32'hff08787f) == 32'h500002b;
wire dec_aesmix_dec  = (encoded & 32'hff08787f) == 32'h508002b;
wire dec_ldr_bu      = (encoded & 32'h3e00787f) == 32'h200002b;
wire dec_ldr_hu      = (encoded & 32'h3e00787f) == 32'h1200002b;
wire dec_ldr_w       = (encoded & 32'hfe00787f) == 32'h2200002b;
wire dec_str_b       = (encoded & 32'h3e00787f) == 32'h200082b;
wire dec_str_h       = (encoded & 32'h3e00787f) == 32'h1200082b;
wire dec_str_w       = (encoded & 32'hfe00787f) == 32'h2200082b;
wire dec_scatter_b   = (encoded & 32'hff00787f) == 32'ha00082b;
wire dec_gather_b    = (encoded & 32'hff00787f) == 32'ha00002b;
wire dec_scatter_h   = (encoded & 32'hff00787f) == 32'hb00082b;
wire dec_gather_h    = (encoded & 32'hff00787f) == 32'hb00002b;
wire dec_bop         = (encoded & 32'h8787f) == 32'h682b;
wire dec_mequ        = (encoded & 32'hf000707f) == 32'h702b;
wire dec_mlte        = (encoded & 32'hf000707f) == 32'h1000702b;
wire dec_mgte        = (encoded & 32'hf000707f) == 32'h2000702b;
wire dec_lut         = (encoded & 32'hf008787f) == 32'h3008702b;
wire dec_madd_3      = (encoded & 32'hf0087c7f) == 32'h4000702b;
wire dec_msub_3      = (encoded & 32'hf0087c7f) == 32'h6000702b;
wire dec_madd_2      = (encoded & 32'hff087c7f) == 32'h5000702b;
wire dec_msub_2      = (encoded & 32'hff087c7f) == 32'h5100702b;
wire dec_macc_2      = (encoded & 32'hff087c7f) == 32'h5200702b;
wire dec_macc_1      = (encoded & 32'hfff87c7f) == 32'h5f00702b;
wire dec_msll        = (encoded & 32'hf0087c7f) == 32'h7000782b;
wire dec_msrl        = (encoded & 32'hf0087c7f) == 32'h8000782b;
wire dec_mmul_3      = (encoded & 32'hf0087c7f) == 32'h9000782b;
wire dec_mclmul_3    = (encoded & 32'hf0087c7f) == 32'ha000782b;
wire dec_msll_i      = (encoded & 32'hc0087c7f) == 32'hc000742b;
wire dec_msrl_i      = (encoded & 32'hc0087c7f) == 32'h8000742b;
wire dec_ld_bu       = (encoded & 32'h707f) == 32'h102b;
wire dec_ld_hu       = (encoded & 32'h10707f) == 32'h202b;
wire dec_ld_w        = (encoded & 32'h10787f) == 32'h302b;
wire dec_ld_hiu      = (encoded & 32'h10787f) == 32'h10302b;
wire dec_ld_liu      = (encoded & 32'h10787f) == 32'h10382b;
wire dec_ipbit       = (encoded & 32'h7f8787f) == 32'h10202b;
wire dec_pbit        = (encoded & 32'h7f8787f) == 32'h10282b;
wire dec_pbyte       = (encoded & 32'hf8787f) == 32'h30202b;
wire dec_ins         = (encoded & 32'h38787f) == 32'h30282b;
wire dec_bmv         = (encoded & 32'h38787f) == 32'h38202b;
wire dec_ext         = (encoded & 32'h38787f) == 32'h38282b;
wire dec_st_b        = (encoded & 32'h707f) == 32'h402b;
wire dec_st_h        = (encoded & 32'h100707f) == 32'h502b;
wire dec_st_w        = (encoded & 32'h100787f) == 32'h602b;
wire [3:0] dec_arg_crs3    = encoded[27:24];
wire [2:0] dec_arg_pw      = encoded[31:29];
wire [3:0] dec_arg_crs1    = encoded[18:15];
wire [7:0] dec_arg_lut8    = encoded[31:24];
wire [1:0] dec_arg_b0      = encoded[31:30];
wire [3:0] dec_arg_crd     = encoded[10:7];
wire [4:0] dec_arg_imm5    = encoded[19:15];
wire [5:0] dec_arg_cmshamt = encoded[29:24];
wire [4:0] dec_arg_rd      = encoded[11:7];
wire [2:0] dec_arg_crdm    = encoded[9:7];
wire [4:0] dec_arg_cl      = encoded[26:22];
wire [1:0] dec_arg_b2      = encoded[27:26];
wire [4:0] dec_arg_rs1     = encoded[19:15];
wire [0:0] dec_arg_cc      = encoded[11:11];
wire [3:0] dec_arg_crs2    = encoded[23:20];
wire [4:0] dec_arg_cshamt  = encoded[24:20];
wire [1:0] dec_arg_b3      = encoded[25:24];
wire [4:0] dec_arg_rs2     = encoded[24:20];
wire [10:0] dec_arg_imm11   = encoded[31:21];
wire [0:0] dec_arg_ca      = encoded[24:24];
wire [3:0] dec_arg_imm11lo = encoded[10:7];
wire [4:0] dec_arg_cs      = encoded[31:27];
wire [6:0] dec_arg_imm11hi = encoded[31:25];
wire [0:0] dec_arg_cd      = encoded[20:20];
wire [1:0] dec_arg_b1      = encoded[29:28];
wire dec_invalid_opcode = !(dec_bop || dec_msrl || dec_padd || dec_aessub_encrot || dec_msub_3 || dec_madd_2 || dec_sha3_xy || dec_psrl || dec_psll_i || dec_gpr2xcr || dec_ins || dec_ld_w || dec_prot || dec_str_h || dec_rngsamp || dec_ldr_bu || dec_ld_bu || dec_ld_hiu || dec_ext || dec_ldr_hu || dec_sha3_x2 || dec_madd_3 || dec_pbit || dec_msrl_i || dec_st_b || dec_pmul_l || dec_rngseed || dec_psll || dec_rngtest || dec_macc_1 || dec_sha3_x4 || dec_init || dec_aessub_enc || dec_bmv || dec_xcr2gpr || dec_aessub_dec || dec_str_b || dec_mclmul_3 || dec_sha3_x1 || dec_pmul_h || dec_mmul_3 || dec_msll_i || dec_aesmix_enc || dec_gather_b || dec_ld_liu || dec_scatter_b || dec_ipbit || dec_mequ || dec_pclmul_h || dec_mgte || dec_pclmul_l || dec_sha3_yx || dec_cmov_f || dec_psub || dec_msub_2 || dec_msll || dec_ld_hu || dec_aessub_decrot || dec_aesmix_dec || dec_macc_2 || dec_st_h || dec_pbyte || dec_gather_h || dec_lut || dec_st_w || dec_prot_i || dec_psrl_i || dec_cmov_t || dec_scatter_h || dec_str_w || dec_mlte || dec_ldr_w);
